`define  FORMAL  1
`define  COREV_ASSERT_OFF  1 // TEMP: To avoid errors, only chech reference model assertions
`define  QUESTA_VSIM 1 // Also solves problems with onespin